localparam NUM_COMPARISONS = 256;
localparam NUM_ROTATIONS = 64;
localparam bit signed [4:0] ORB_SAMPLES [NUM_COMPARISONS][2][2] = '{
	'{'{3,8},'{-5,9}},
	'{'{-2,4},'{12,7}},
	'{'{-9,-11},'{-2,-8}},
	'{'{12,7},'{13,12}},
	'{'{13,2},'{-12,2}},
	'{'{7,1},'{-6,1}},
	'{'{10,-2},'{4,-2}},
	'{'{13,-13},'{8,-11}},
	'{'{3,-13},'{9,-12}},
	'{'{-4,10},'{-9,11}},
	'{'{8,-13},'{9,-8}},
	'{'{-7,-11},'{-12,-9}},
	'{'{-7,7},'{-6,12}},
	'{'{5,-4},'{0,-3}},
	'{'{-2,-13},'{3,-12}},
	'{'{0,-9},'{-5,-7}},
	'{'{6,12},'{1,12}},
	'{'{-6,-3},'{-12,-2}},
	'{'{13,-6},'{8,-4}},
	'{'{13,11},'{8,12}},
	'{'{-7,4},'{-1,5}},
	'{'{3,5},'{3,10}},
	'{'{7,3},'{-12,6}},
	'{'{7,-8},'{2,-6}},
	'{'{-11,-2},'{10,-1}},
	'{'{-12,-13},'{-10,-8}},
	'{'{-3,-7},'{3,-5}},
	'{'{-2,-4},'{-7,-3}},
	'{'{12,-10},'{-11,-6}},
	'{'{12,5},'{7,6}},
	'{'{6,5},'{1,7}},
	'{'{0,1},'{5,4}},
	'{'{-11,9},'{13,11}},
	'{'{-7,4},'{-12,4}},
	'{'{1,2},'{-4,4}},
	'{'{12,-4},'{-7,-2}},
	'{'{5,-8},'{10,-7}},
	'{'{-11,4},'{-12,9}},
	'{'{8,0},'{13,1}},
	'{'{2,-13},'{-2,-8}},
	'{'{2,-3},'{-3,-2}},
	'{'{-9,-6},'{9,-4}},
	'{'{-12,8},'{-7,10}},
	'{'{-9,0},'{-3,1}},
	'{'{5,7},'{10,11}},
	'{'{6,-13},'{0,-11}},
	'{'{-7,10},'{-1,12}},
	'{'{3,-6},'{-12,-6}},
	'{'{9,10},'{4,12}},
	'{'{-8,-13},'{12,-8}},
	'{'{0,-13},'{4,-8}},
	'{'{-3,3},'{-8,7}},
	'{'{-7,5},'{7,10}},
	'{'{-7,-1},'{12,1}},
	'{'{10,3},'{-6,5}},
	'{'{4,2},'{10,3}},
	'{'{0,-13},'{-5,-13}},
	'{'{7,-13},'{-12,-12}},
	'{'{-3,-13},'{-8,-11}},
	'{'{-12,-7},'{-7,-4}},
	'{'{10,6},'{-8,12}},
	'{'{1,-9},'{6,-7}},
	'{'{5,-2},'{-12,0}},
	'{'{-5,-12},'{-5,-7}},
	'{'{10,3},'{13,8}},
	'{'{7,-7},'{-5,-4}},
	'{'{2,-3},'{7,-1}},
	'{'{-9,2},'{11,5}},
	'{'{13,-11},'{13,-5}},
	'{'{-6,-1},'{1,0}},
	'{'{3,5},'{-2,5}},
	'{'{13,-4},'{-12,-4}},
	'{'{6,-9},'{-6,-9}},
	'{'{10,-12},'{4,-8}},
	'{'{-2,10},'{3,12}},
	'{'{-12,7},'{-12,12}},
	'{'{13,-7},'{-5,-6}},
	'{'{-9,-4},'{-4,-3}},
	'{'{1,7},'{-2,12}},
	'{'{-6,-7},'{-1,-5}},
	'{'{-11,-13},'{-5,-12}},
	'{'{-7,-3},'{6,-2}},
	'{'{8,7},'{7,12}},
	'{'{7,-13},'{12,-11}},
	'{'{3,1},'{-12,12}},
	'{'{6,2},'{0,3}},
	'{'{-3,-4},'{13,-2}},
	'{'{13,-1},'{-9,1}},
	'{'{-1,7},'{6,8}},
	'{'{1,1},'{-12,3}},
	'{'{-1,9},'{-6,12}},
	'{'{9,-1},'{-3,-1}},
	'{'{13,-13},'{-5,-10}},
	'{'{-7,7},'{-12,10}},
	'{'{5,12},'{-9,12}},
	'{'{-3,6},'{-11,7}},
	'{'{13,5},'{-10,6}},
	'{'{12,2},'{-3,2}},
	'{'{-8,3},'{6,4}},
	'{'{-6,2},'{13,12}},
	'{'{12,9},'{-3,10}},
	'{'{-4,-8},'{-9,-7}},
	'{'{-12,-11},'{6,-4}},
	'{'{-12,1},'{8,2}},
	'{'{9,6},'{4,7}},
	'{'{-3,2},'{2,3}},
	'{'{-3,6},'{0,11}},
	'{'{3,3},'{8,8}},
	'{'{-8,7},'{-3,9}},
	'{'{5,-11},'{4,-6}},
	'{'{-11,-10},'{-10,-5}},
	'{'{8,-5},'{-12,-3}},
	'{'{-5,-10},'{0,-9}},
	'{'{1,8},'{6,12}},
	'{'{6,4},'{11,6}},
	'{'{-12,-10},'{-7,-8}},
	'{'{2,4},'{-7,6}},
	'{'{0,-2},'{-12,-2}},
	'{'{8,-5},'{-2,-5}},
	'{'{6,7},'{-12,10}},
	'{'{13,-9},'{8,-8}},
	'{'{13,-5},'{2,-5}},
	'{'{8,8},'{13,9}},
	'{'{11,-9},'{0,-9}},
	'{'{8,1},'{2,1}},
	'{'{4,7},'{-1,9}},
	'{'{-1,-2},'{4,-1}},
	'{'{6,11},'{11,12}},
	'{'{9,-12},'{-4,-6}},
	'{'{-7,3},'{-12,7}},
	'{'{-5,5},'{-8,10}},
	'{'{4,0},'{-8,2}},
	'{'{-12,-9},'{13,-5}},
	'{'{-7,0},'{-12,2}},
	'{'{-2,-1},'{-7,1}},
	'{'{-11,5},'{9,7}},
	'{'{-5,3},'{8,6}},
	'{'{4,-13},'{-9,-8}},
	'{'{-9,-5},'{3,-3}},
	'{'{7,-4},'{12,-3}},
	'{'{-5,6},'{0,8}},
	'{'{-6,-7},'{-12,-6}},
	'{'{-6,-13},'{2,-5}},
	'{'{10,1},'{-10,3}},
	'{'{-1,4},'{4,8}},
	'{'{2,-2},'{13,2}},
	'{'{12,2},'{-12,12}},
	'{'{13,-2},'{6,0}},
	'{'{-1,4},'{-3,9}},
	'{'{10,-6},'{5,-3}},
	'{'{13,-3},'{-1,-1}},
	'{'{-5,7},'{11,12}},
	'{'{2,4},'{7,5}},
	'{'{-9,-13},'{5,-9}},
	'{'{-1,7},'{-6,8}},
	'{'{8,7},'{-6,7}},
	'{'{4,-7},'{-1,-7}},
	'{'{-11,-8},'{8,-7}},
	'{'{-6,-13},'{8,-12}},
	'{'{-4,2},'{-9,3}},
	'{'{5,10},'{-3,12}},
	'{'{5,-6},'{-7,-6}},
	'{'{3,8},'{8,9}},
	'{'{12,2},'{-8,2}},
	'{'{2,-11},'{-3,-10}},
	'{'{13,-12},'{9,-7}},
	'{'{0,-11},'{5,-10}},
	'{'{3,5},'{-8,11}},
	'{'{13,-2},'{-12,-1}},
	'{'{8,-1},'{-9,0}},
	'{'{11,-13},'{5,-12}},
	'{'{2,-10},'{-11,-10}},
	'{'{-9,-3},'{13,-2}},
	'{'{3,2},'{-2,3}},
	'{'{13,-9},'{0,-4}},
	'{'{-6,-4},'{10,-3}},
	'{'{-12,-4},'{7,-2}},
	'{'{11,-6},'{-9,-4}},
	'{'{3,6},'{-11,6}},
	'{'{-11,-13},'{-5,-5}},
	'{'{-11,11},'{-6,12}},
	'{'{5,7},'{2,12}},
	'{'{-12,-1},'{-7,0}},
	'{'{8,-4},'{2,-3}},
	'{'{-1,-7},'{-7,-6}},
	'{'{12,-13},'{13,-8}},
	'{'{2,-7},'{8,-6}},
	'{'{-5,-8},'{9,-6}},
	'{'{1,-5},'{-5,-4}},
	'{'{-7,-13},'{-10,-8}},
	'{'{-5,1},'{13,5}},
	'{'{0,1},'{13,10}},
	'{'{-12,9},'{1,10}},
	'{'{8,5},'{9,10}},
	'{'{-11,-1},'{13,1}},
	'{'{3,-9},'{-2,-6}},
	'{'{10,-1},'{-12,1}},
	'{'{-1,-13},'{10,-8}},
	'{'{11,8},'{6,10}},
	'{'{13,2},'{6,3}},
	'{'{13,7},'{9,12}},
	'{'{10,-10},'{7,-5}},
	'{'{8,-10},'{13,-8}},
	'{'{6,4},'{-5,8}},
	'{'{-12,3},'{13,8}},
	'{'{-2,-4},'{3,-3}},
	'{'{13,5},'{12,10}},
	'{'{13,4},'{1,5}},
	'{'{-9,-9},'{-3,-4}},
	'{'{-3,0},'{9,3}},
	'{'{-1,-12},'{-1,-6}},
	'{'{-2,3},'{8,4}},
	'{'{10,-10},'{-9,-10}},
	'{'{13,8},'{-12,12}},
	'{'{12,-8},'{5,-6}},
	'{'{-2,2},'{-7,3}},
	'{'{-6,10},'{8,11}},
	'{'{-8,6},'{12,8}},
	'{'{-10,-7},'{-5,-6}},
	'{'{9,-3},'{-9,-3}},
	'{'{13,-1},'{-5,-1}},
	'{'{7,-3},'{-4,-3}},
	'{'{2,-8},'{-3,-8}},
	'{'{-2,4},'{-12,12}},
	'{'{5,2},'{-11,3}},
	'{'{9,6},'{13,11}},
	'{'{1,3},'{-12,7}},
	'{'{1,11},'{-4,12}},
	'{'{0,-3},'{-6,-3}},
	'{'{11,4},'{-12,4}},
	'{'{4,2},'{-1,2}},
	'{'{6,-10},'{-1,-8}},
	'{'{-7,-13},'{-1,-11}},
	'{'{-12,-13},'{13,-11}},
	'{'{0,6},'{13,11}},
	'{'{1,0},'{-4,1}},
	'{'{-3,-13},'{2,-9}},
	'{'{-8,-9},'{3,-6}},
	'{'{6,-13},'{2,-8}},
	'{'{9,5},'{-10,8}},
	'{'{-7,2},'{9,3}},
	'{'{6,-1},'{1,-1}},
	'{'{-5,9},'{2,11}},
	'{'{3,11},'{8,12}},
	'{'{0,3},'{-5,3}},
	'{'{-4,-1},'{-10,0}},
	'{'{6,3},'{-5,4}},
	'{'{0,-13},'{-5,-10}},
	'{'{-8,5},'{-11,12}},
	'{'{-9,8},'{6,9}},
	'{'{4,7},'{12,8}},
	'{'{-4,-10},'{-9,-10}},
	'{'{-3,7},'{-4,12}},
	'{'{7,9},'{2,10}},
	'{'{0,7},'{2,12}},
	'{'{6,-1},'{1,0}}
};

localparam bit signed [8:0] ROTATION_LUT [NUM_ROTATIONS][2] = '{
	'{255,0},
	'{255,25},
	'{251,50},
	'{245,74},
	'{237,98},
	'{226,121},
	'{213,142},
	'{198,162},
	'{181,181},
	'{162,198},
	'{142,213},
	'{121,226},
	'{98,237},
	'{74,245},
	'{50,251},
	'{25,255},
	'{0,255},
	'{-25,255},
	'{-50,251},
	'{-74,245},
	'{-98,237},
	'{-121,226},
	'{-142,213},
	'{-162,198},
	'{-181,181},
	'{-198,162},
	'{-213,142},
	'{-226,121},
	'{-237,98},
	'{-245,74},
	'{-251,50},
	'{-255,25},
	'{-256,0},
	'{-255,-25},
	'{-251,-50},
	'{-245,-74},
	'{-237,-98},
	'{-226,-121},
	'{-213,-142},
	'{-198,-162},
	'{-181,-181},
	'{-162,-198},
	'{-142,-213},
	'{-121,-226},
	'{-98,-237},
	'{-74,-245},
	'{-50,-251},
	'{-25,-255},
	'{0,-256},
	'{25,-255},
	'{50,-251},
	'{74,-245},
	'{98,-237},
	'{121,-226},
	'{142,-213},
	'{162,-198},
	'{181,-181},
	'{198,-162},
	'{213,-142},
	'{226,-121},
	'{237,-98},
	'{245,-74},
	'{251,-50},
	'{255,-25}
};
